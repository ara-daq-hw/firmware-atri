`timescale 1ns / 1ps
// sigh attempt to make a trigger that actually works?
module trigger_scaler_v3(
		input trigger_i,
		input power_i,
		input mask_i,
		output trig_p_o,
		output trig_n_o,
		output scaler_o,
		
		input fast_clk_i,
		input slow_clk_i,
		input slow_ce_i,
		// This is unused. It's here for compatibility with trigger_scaler_v4.
		input trig_oneshot_i
    );
	 
	// Bleah, this is crap. Just do this the sleazy way. Self-disabling latch, that gets synchronized
	// and then cleared. The synchronized copy starts a shift register. If a new trigger occurs, reset
	// the shreg. If the shreg reaches 3 cycles, reset the shreg.
	// Trigger is generated by a latch that self-disables.

	wire trig_bit;
	wire trig_clr;
	LDCE #(.INIT(0)) trig_latch(.D(trigger_i),.GE(power_i),.G(!trig_bit),.Q(trig_bit),.CLR(trig_clr));
	parameter ONE_SHOT_LENGTH = 3;
	reg [1:0] trig_sync = {2{1'b0}};
	reg [ONE_SHOT_LENGTH-1:0] trig_shreg = {ONE_SHOT_LENGTH{1'b0}};
	reg trigger_output = 0;

	always @(posedge fast_clk_i) begin
		if (trig_sync[1:0] == 2'b01) trig_sync[1] <= 1;
		else trig_sync[1] <= 0;
		trig_sync <= {trig_sync[0],trig_bit};
	end
	assign trig_clr = trig_sync[1];
	// Set the beginning bit if we see a trigger. ONLY clear it if we see the top bit of the
	// shreg go.
	always @(posedge fast_clk_i) begin
		if (trig_sync[1]) trigger_output <= 1;
		else if (trig_shreg[ONE_SHOT_LENGTH-1]) trigger_output <= 0;
	end
	always @(posedge fast_clk_i) begin
		if (trig_shreg[ONE_SHOT_LENGTH-1] || trig_sync[1])
			trig_shreg[ONE_SHOT_LENGTH-1:0] <= {ONE_SHOT_LENGTH{1'b0}};
		else
			trig_shreg <= {trig_shreg[ONE_SHOT_LENGTH-2:0],trigger_output};
	end
	//% Indicates that the flag is still traversing the synchronizer.
	wire busy_p;
	//% Flags in the slow clock domain for the +/- edge clear flags. Both on +edge of slowclk.
	wire p_cleared_slowclk;
	//% Flag generator to inform slow clock that positive edge chain has seen a clear.
	flag_sync clear_p_flag(.clkA(fast_clk_i),.clkB(slow_clk_i),.in_clkA(trig_shreg[ONE_SHOT_LENGTH-1] && !busy_p),
									.out_clkB(p_cleared_slowclk),.busy_clkA(busy_p));

	//% Generates a scaler output, with stuck-on detection. No higher level trigger needs this.
	scaler_generator sc_gen(.trig_i(trigger_output),
									.fclk_i(fast_clk_i),.sclk_i(slow_clk_i),
									.sce_i(slow_ce_i),
									.clear_sclk_i(p_cleared_slowclk),
									.scaler_o(scaler_o));

	assign trig_p_o = trigger_output;
endmodule
