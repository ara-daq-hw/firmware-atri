`define EVIF_SIZE 63
