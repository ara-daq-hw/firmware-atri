`timescale 1ns / 1ps
`include "trigger_defs.vh"
// Trigger_scaler_v5.
// v5 adds per-channel trigger delay value inputs.
module trigger_scaler_v5(
		trigger_i,
		power_i,
		mask_i,
		trig_p_o,
		trig_n_o,
		scaler_o,
		
		fast_clk_i,
		slow_clk_i,
		slow_ce_i,
		sync_i,
		delay_i,
		trig_oneshot_i
    );
	parameter ONE_SHOT_MAX_BITS = `TRIG_ONESHOT_BITS;
	parameter TRIG_DELAY_VAL_BITS = `TRIG_DELAY_VAL_BITS;
	parameter POLARITY = "POSITIVE";
	
	input trigger_i;
	input power_i;
	input mask_i;
	output trig_p_o;
	output trig_n_o;
	output scaler_o;
	
	input fast_clk_i;
	input slow_clk_i;
	input slow_ce_i;
	input sync_i;
	input [TRIG_DELAY_VAL_BITS-1:0] delay_i;
	input [ONE_SHOT_MAX_BITS-1:0] trig_oneshot_i;
	
	// Bleah, this is crap. Just do this the sleazy way. Self-disabling latch, that gets synchronized
	// and then cleared. The synchronized copy starts a shift register. If a new trigger occurs, reset
	// the shreg. If the shreg reaches 3 cycles, reset the shreg.
	// Trigger is generated by a latch that self-disables.

	///// POSITIVE POLARITY
	wire trig_bit;
	wire trig_reset;
	reg [1:0] trig_sync = {2{1'b0}};
	reg [ONE_SHOT_MAX_BITS-1:0] trig_count = {ONE_SHOT_MAX_BITS{1'b0}};
	(* EQUIVALENT_REGISTER_REMOVAL = "NO" *)
	reg [ONE_SHOT_MAX_BITS-1:0] trig_oneshot_sync = {ONE_SHOT_MAX_BITS{1'b0}};
	reg trigger_output = 0;
	reg trigger_unmasked = 0;
	wire trig_valid;
	generate
		if (POLARITY == "POSITIVE") begin : POS
			(* IOB = "TRUE" *)
			LDCE #(.INIT(0)) trig_latch(.D(trigger_i),.GE(power_i),.G(!trig_bit),.Q(trig_bit),.CLR(trig_reset));
			// Synchronize the input trigger. We probably
			// need to add a second synchronizer stage here...
			always @(posedge fast_clk_i) begin
				if (trig_sync[1:0] == 2'b01) trig_sync[1] <= 1;
				else trig_sync[1] <= 0;
				trig_sync[0] <= trig_bit;
			end
			assign trig_reset = trig_sync[1];
			assign trig_valid = trig_sync[1] && power_i;
		end else begin : NEG
			(* IOB = "TRUE" *)
			LDPE #(.INIT(1)) trig_latch(.D(trigger_i),.GE(power_i),.G(trig_bit),.Q(trig_bit),.PRE(trig_reset));
			// Synchronize the input trigger. We probably need to
			// add a second synchronizer stage here...
			always @(posedge fast_clk_i) begin
				if (trig_sync[1:0] == 2'b00) trig_sync[1] <= 1;
				else trig_sync[1] <= 0;
				trig_sync[0] <= trig_bit;
			end
			assign trig_reset = trig_sync[1];
			assign trig_valid = trig_sync[1] && power_i;
		end
	endgenerate
	
	// Synchronize the number of bits we're supposed to wait.
	always @(posedge fast_clk_i) begin
		trig_oneshot_sync <= trig_oneshot_i;
	end

	// Set the beginning bit if we see a trigger. ONLY clear it if we see the top bit of the
	// shreg go, or if the mask turns on.
	always @(posedge fast_clk_i) begin
		if (trig_valid && !mask_i) trigger_output <= 1;
		else if ((trig_count == trig_oneshot_sync) || (mask_i)) trigger_output <= 0;
	end
	// Copy of trigger_output, but non-masked.
	always @(posedge fast_clk_i) begin
		if (trig_valid) trigger_unmasked <= 1;
		else if (trig_count == trig_oneshot_sync) trigger_unmasked <= 0;
	end
	
	// This is the clear for the *unmasked* trigger.
	always @(posedge fast_clk_i) begin
		if ((trig_count == trig_oneshot_sync) || (trig_valid))
			trig_count  <= {ONE_SHOT_MAX_BITS{1'b0}};
		else if (trigger_unmasked)
			trig_count <= trig_count + 1;
	end

	//% Indicates that the flag is still traversing the synchronizer.
	wire busy_p;
	//% Flags in the slow clock domain for the +/- edge clear flags. Both on +edge of slowclk.
	wire p_cleared_slowclk;
	//% Delayed trigger.
	wire trigger_delayed;

	SRLC32E #(.INIT(32'h00000000)) trigger_delay(.D(trigger_output),
																.A(delay_i),
																.CLK(fast_clk_i),
																.Q(trigger_delayed));																

	//% Flag generator to inform slow clock that positive edge chain has seen a clear.
	flag_sync clear_p_flag(.clkA(fast_clk_i),.clkB(slow_clk_i),.in_clkA(trig_count == trig_oneshot_sync && !busy_p),
									.out_clkB(p_cleared_slowclk),.busy_clkA(busy_p));

	//% Generates a scaler output, with stuck-on detection. No higher level trigger needs this.
	scaler_generator sc_gen(.trig_i(trigger_unmasked),
									.fclk_i(fast_clk_i),.sclk_i(slow_clk_i),
									.sce_i(slow_ce_i),
									.sync_i(sync_i),
									.clear_sclk_i(p_cleared_slowclk),
									.scaler_o(scaler_o));

	assign trig_p_o = trigger_delayed;
endmodule
