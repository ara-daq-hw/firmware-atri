`define I2CIF_SIZE 21
