
		.INIT_00(256'h401450A62001401054064001601F501620014005C001C0000001500020204000),
		.INIT_01(256'h46060112000A0401030002CB0104E01540044604400654CD2010401550062001),
		.INIT_02(256'h011200080400030102030140C018000001250006400650614611503C46015026),
		.INIT_03(256'h46040104C001601540060176011D0203011200000112000A01CB0112000A0130),
		.INIT_04(256'h8008410440044004C003C0030000013B61150001012500004006012150444608),
		.INIT_05(256'h01761919C11A6115020300000112C00460150400030002030104C103C003A100),
		.INIT_06(256'h43595075435840060121506D421B43044204420442040104E015C00460154006),
		.INIT_07(256'h0000152140006015010401120401030102C001CB000A4006012150A3435A5093),
		.INIT_08(256'h0176011204000301020301400020C0180020016A01200058013B012800110125),
		.INIT_09(256'h4011C011C012C004601501210004500611214200621F010460154006E01F0001),
		.INIT_0A(256'h4180E0184080E0174080E016408001250000017F4006012160154006509F2001),
		.INIT_0B(256'hC0056015C0036018C0036017C0036016016A61150059013B00118108E1158105),
		.INIT_0C(256'h0000017FC014400601761919C1126115C003408001120400030002030180C003),
		.INIT_0D(256'h00DEE223E122621A6119E01B800111084000E021601BE020C040A00F40150125),
		.INIT_0E(256'h013B00111100800CE015E21AE119E200D100E21B1010A20091005CE9E200D100),
		.INIT_0F(256'hC203521001816015C0036023C0036022C0036021C0036020016A81046115005A),
		.INIT_10(256'hC1206120E21AE1190200010642834181400601761919C10E611554FEC001E102),
		.INIT_11(256'h551DC101D0208101E1FF000002034112B000C00192409130D5205510A000E120),
		.INIT_12(256'h0301020301CBC00100D5011D0201010700550185E01CA0005521C0015210A000),
		.INIT_13(256'h413B403AE11D8114E01CA000C003601CC0030008011200060130011200060400),
		.INIT_14(256'hC2030245E000F130F02063116212F130F02063136214E100F020621DD020621C),
		.INIT_15(256'hC003C103C203621CC2030280C203C203C203C2030200C203621DC203C2030200),
		.INIT_16(256'hC003C203C003C203021B8108A0000112000401D1011200040400030102030136),
		.INIT_17(256'h000AA000C0000041011200040400030002010121A000C003C003C103C0030000),
		.INIT_18(256'h0000000000000000000000000000A00051852010400041120401030102CB01C0),
		.INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_30(256'h4901577D49014901577D49004901530629014902437D532E4900530649064924),
		.INIT_31(256'h036C0D010C000BF00A01090A577D4901490103680903577D49004901577D4908),
		.INIT_32(256'h29024902437D036CC904090A0D000C010B040AF0C9040906577D037303680906),
		.INIT_33(256'hE93A537D5B7DC9144901577D490049014901577D49454901537D49014925532E),
		.INIT_34(256'h036C09040D010C000BF60A0149014901437D53484F0153484F114F0103680905),
		.INIT_35(256'h0B040AF6036C09060D000C010B040A28CF046F3ACF04535229084900577D0373),
		.INIT_36(256'h9BD09AC0DEB05EA04368B000C9014A01437D036C693A0C000B040A01036C0904),
		.INIT_37(256'h8001C900090343758A01B000CB01B40059C05CA049010A360B04436CB000C901),
		.INIT_38(256'h0000000000000000000000000000000000000000000000000200040600080100),
		.INIT_39(256'h00000000000000000000004B4F20302E31762050445520657A616C426F636950),
		.INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_3F(256'h4300000000000000000000000000000000000000000000000000000000000000),
		.INITP_00(256'h343003F777F40093F40D002940A30CFD04FC0C30C008CF7770020F4D34D34E34),
		.INITP_01(256'h808888D0C1A96175282762033BF48C024888C31922233F3D2933D038F00230C3),
		.INITP_02(256'h28C00AA8AA1B0C00A88AA2288541414409A88C3002303AD2D903958A0AA0FD34),
		.INITP_03(256'h000000000000000000000000000000000000000000000000000000000002D300),
		.INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INITP_06(256'hE366403958E4F00C0C008B4FC000F74CBD3434D34F8008FCC00D334D34D34F74),
		.INITP_07(256'hC000000000000000000000000000000000000000000000000000000000000000)		