
		.INIT_00(256'h50122002400154082001400950144C204D43CC430C00090008000B000A000E00),
		.INIT_01(256'hF200D3104350425101FFC03F000C000CC001101000DF404240F100FF40080026),
		.INIT_02(256'h503084015C34020E04000310424200C30F000E454008CC430C00400858235023),
		.INIT_03(256'h010600DF6002AA009A400A080B0E0A080B0E542C431483019B10F13000DFE0FF),
		.INIT_04(256'h4050544C20014024505D4E455457200240015457200140098B008A04AB009A10),
		.INIT_05(256'h404CAB008A05405D0E4F404C0E46505B4E45404CCC430C205C62F1B0D0A04151),
		.INIT_06(256'hC081C180010250804E4650804E42CB81CA80EB00CA02CE81C08010F000F100FE),
		.INIT_07(256'hA8008801C981C880C1816106C1806105C1816108C1806107C1816104C1806103),
		.INIT_08(256'hC3814367C3804366C2605C94010E820102FFB1D0C1816102C180010E010E6101),
		.INIT_09(256'h50A22202C181D1C0D12002064242A1016101C18061005488C3814365C3804364),
		.INIT_0A(256'hE0206000C023601350AE2210C022601250AA2208C021601150A62204C0206010),
		.INIT_0B(256'hB0004E4FB0004E4654B85010414040420B000A00C0240001C001E021A0016001),
		.INIT_0C(256'hE0024002E0014001E0004000C14110FF4E455460F0104142404040280E428F01),
		.INIT_0D(256'h0100A000C0090002E0084008E0074007E0064006E0054005E0044004E0034003),
		.INIT_0E(256'hA100000EA100000EA100000EA100000EA100000EA100000EA100000EA100000E),
		.INIT_0F(256'h407040FEC181C082C1810100C1800101C1810100C180015858F141034150A000),
		.INIT_10(256'h000000000000000000000000000000008000C7316721C7306720A0005500C001),
		.INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_3F(256'h410340F100FD0000000000000000000000000000000000000000000000000000),
		.INITP_00(256'h5A888888A376968CD73378D434DD3455B16AB56C1E030E3F500A4CCFD34D2000),
		.INITP_01(256'h3A8888D26666666628888888888B703199D008E088D8D8D8D820238888B908A8),
		.INITP_02(256'h000000000000000000000000000000000000000000000000000000000000E22D),
		.INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INITP_07(256'hF000000000000000000000000000000000000000000000000000000000000000)		