
		.INIT_00(256'h007E14D12002006F007E14AB2004006F402140040007001300D9C001033E0F38),
		.INIT_01(256'h50264000A000001EE00A4080E0094080E0084080B40020014011A00014C82001),
		.INIT_02(256'hE00910A0CA026A09690B404F502B2001E00B408040224E80B000C00160094021),
		.INIT_03(256'h600BC0800000C0800003C0806008544700E55432C0018101F21042800110035B),
		.INIT_04(256'h408040440010C08000FFC0800001C0806008A000C01100104044C0806009C080),
		.INIT_05(256'h6009C080600BC0800000C08080026009C0806008544700E503451A00690BE009),
		.INIT_06(256'hF0F08F01F1F08F01F2F08F01F3F040445463C0018101C280721001105044C000),
		.INIT_07(256'h70F0CF01A00071F0CF01007EA00072F0CF01007AA00073F0CF010076A0008F01),
		.INIT_08(256'hB020913040898401588EF020D1300400A0009010408282015886D0100200A000),
		.INIT_09(256'h6E00A000EE00BE006E00A000000E000E000E000EA0000006000600060006A000),
		.INIT_0A(256'hE0100030035B0A02091CA00000E5E0100001E011035B0A020982A000EE00DE00),
		.INIT_0B(256'hE0100003035B0A02098200A3E10C0101000540B90100000450B700E5E0110000),
		.INIT_0C(256'h54C600A3000400A30005B0004001600C409B00F7409F000854C600E5E0110000),
		.INIT_0D(256'hE011000FE0100039035B0A0209C040C454C600A3C004600C00A3C006600C40C4),
		.INIT_0E(256'h00000000000000000000000000000000A00058E54801A000C020000458E04801),
		.INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INIT_32(256'hA000C8040890C903000000000000000000000000000000000000000000000000),
		.INIT_33(256'hC8010800A000C8040840A000C804C84057390810C803A000C804C84857330820),
		.INIT_34(256'h03305B794A01577028A0A00008000910C838084B032CA000C80208C0C8000818),
		.INIT_35(256'h08000910C8380861032C434DCA018901F89048035770282080010800C8380854),
		.INIT_36(256'h43618901CA01577028A080010800C838086B033578905B794A01577028A0A000),
		.INIT_37(256'h437D4804800180010801C838087280010800C8380872033B8001080257744A01),
		.INIT_38(256'h000000000000000000000000000000000000000000737365726464412043414D),
		.INIT_39(256'h000000002E0000002E0000002E00000000000000000073736572646441205049),
		.INIT_3A(256'h000000203A64657265776F5020414444000000203A746E657365725020414444),
		.INIT_3B(256'h000000416D20000000203A4920414444000000562000002E00203A5620414444),
		.INIT_3C(256'h000000203A7365636976654420414444000000432000000000203A5420414444),
		.INIT_3D(256'h00000000000000203A7374656B6361500000000000203A64657463656E6E6F43),
		.INIT_3E(256'h000000002E0000002E0000002E00000000000073736572646441205049204350),
		.INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INITP_00(256'h18787879999BD60D22248FC2322228E22223F583843D8C93DB88892DF7F73FFC),
		.INITP_01(256'h000000000000B68D88C3F0C3F324CCF88C3830F88C2E2C28282AAAAA5DD49DD2),
		.INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.INITP_06(256'hCF2323CDD772337608F58DC8F7608E888A28CA8CA20000000000000000000000),
		.INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000)		