// IRS write controller.

//% @brief IRS write controller.
//%
//% @gensymbol
//% MODULE irs_write_controller_v3
//% LPORT clk_i input
//% LPORT enable_i input
//% LPORT rst_i input
//% LPORT ssp_clk_i input
//% LPORT wrstrb_clk_i input
//% LPORT space
//% LPORT wr_block_i input
//% LPORT wr_phase_o output
//% LPORT wr_ack_o output
//% RPORT ssp_o output
//% RPORT sst_o output
//% RPORT wrstrb_o output
//% RPORT wr_o output
//% @endgensymbol
//%
//% This module outputs a phase (via wr_phase_o) which indicates whether the top half
//% of the sampling cells are being written to, or the bottom half.
//% It also outputs a wr_ack_o signal which indicates that the block which is presented
//% on wr_block_i has been written to.
//%
//% This, therefore, separates the block *fetch* from the block *write*. The block
//% fetching portions are purely digital. These, however, may need to be tuned for optimal
//% timing.
//%
//% It is possible to use the irs_write_controller to write a single block. The timing
//% diagram for this is:
//% @drawtiming
//% clk_i=0,wr_phase_o=1,wr_block_i=X,enable_i=0,wr_ack_o=0,wrstrb=0,sst=0,wr=X.
//% clk_i=1,sst=1.
//% clk_i=0.
//% clk_i=1,wr_phase_o=0.
//% clk_i=0,enable_i=1,wr_block_i="0x004".
//% clk_i=1,sst=0;wr_block_i=>wr="0x000".
//% clk_i=0.
//% clk_i=1,wr_phase_o=1,wrstrb=1,wr_ack_o=1.
//% clk_i=0;wr_ack_o=>enable_i=0;wr_block_i=X.
//% clk_i=1,sst=1,wrstrb=0.
//% clk_i=0.
//% @enddrawtiming
//%
//% Here "enable_i" is just qualified by the write phase of the block write desired - 
//% with an example block of "0x000" (sample cells 0-63), this is wr_phase_o = 0.
//% enable_i is then disabled by being qualified against !wr_ack_o.
//%
//% The write block must be present by the rising clock edge after wr_phase_o first
//% changes (i.e. the third rising clock edge in the diagram above). This is when the
//% block is clocked onto the WR outputs. wr_ack_o is asserted for only one clock cycle
//% (the same clock cycle that WRSTRB is asserted).
//%
//% Nominally, in the previous version of the IRS3 firmware, "ssp_clk_i" is 180 degrees
//% off from clk_i (i.e. CLK180 in a DCM) and wrstrb_clk_i is 270 degrees off from
//% clk_i (i.e. CLK270 in a DCM).
//%
//% Note that the rising edge is used for ssp_clk_i/wrstrb_clk_i.
//%
//% So the base timing there was (starting from the beginning)
//% at   -5 ns: SSp goes high
//% at    0 ns: SSt goes high
//% at   15 ns: SSp goes low
//% at   20 ns: SSt goes low, WR is asserted to the appropriate block.
//% at 27.5 ns: WRSTRB goes high
//% at   35 ns: SSp goes high
//% at 37.5 ns: WRSTRB goes low
//% at   40 ns: SSt goes high, WR is asserted to the appropriate block.
//% at 47.5 ns: WRSTRB goes high
//% at   55 ns: SSp goes low.
//% at 57.5 ns: WRSTRB goes low.
//% etc.
//%
//% Note that WRSTRB and SSp have relatively short timing paths (5 ns and 7.5 ns respectively).
//% Therefore we:
//% 1: register the SSp enable in the clk domain
//% 2: transfer that to the SSp_clk domain
//% This way the only short timing path is from the registered SSp enable-> OBUF, and P&R can
//% just shove it right beside the IOBUF.
//%
//% The WRSTRB timing and width are controllable outside of this module - the delay from a
//% change in SST to WRSTRB is just the delay from clk_i to wrstrb_clk_i, and the width
//% of WRSTRB is just the delay from wrstrb_clk_i to wrstrbn_clk_i.
//% Note that for architectures without a dual-clock DDR flipflop primitive, WRSTRB's width
//% is generated by using an async clear generated by a half-clock-width pulse, so it may be
//% (very) slightly different than expected.
module irs_write_controller_v3(
		// System interface
		input clk_i,					//% System clock (1/32 sampling speed).
		input enable_i, 				//% Begin writing to the IRS.
		input rst_i,					//% System reset.
		input ssp_clk_i,				//% Clock for the SSp timing strobe. Still 4X SSt, but offset in phase.
		input wrstrb_clk_i,			//% Clock for the write strobe going high. Still 4X SSt, offset in phase.
		
		// Interface to the block manager.
		input [8:0] wr_block_i,		//% Block value to use.
		output wr_phase_o,			//% '1' if we need a block for sample cells 64-128, 0 for 0-63
		output wr_ack_o,				//% Block has been written to.
				
		// Interface to the IRS. Connect straight to the IOBUFs for proper timing.
		output ssp_o,					//% Start timing strobe.
		output sst_o,					//% Stop timing strobe.
		output wrstrb_o,				//% Write strobe.
		output [9:0] wr_o,			//% Write lines.

		// Debug outputs. Equivalent to the IRS outputs, except ssp/wrstrb are in clk_i domain.
		output dbg_ssp_o,				//% Debug start timing strobe.
		output dbg_sst_o,				//% Debug stop timing strobe.
		output dbg_wrstrb_o,			//% Debug write strobe.
		output [9:0] dbg_wr_o,		//% Debug write address.
		output [3:0] dbg_state_o	//% Debug state.
		);
	
	//% Determines how WRSTRB is generated. Can be SPARTAN6, SPARTAN3, VIRTEX2, SPARTAN3A, SPARTAN3E, or other.
	parameter ARCH = "SPARTAN6";

	`include "clogb2.vh"
	// WR is latched at the transition into SAMPLE_LOW_PREP_HIGH and PREP_LOW_SAMPLE_HIGH.
	// That means that wr_phase_o needs to be '1' in TRANSFER_LOW_SAMPLE_HIGH and SAMPLE_LOW_PREP_HIGH,
	// and 0 in SAMPLE_LOW_TRANSFER_HIGH and PREP_LOW_SAMPLE_HIGH.
	// wr_phase_o is only high in SAMPLE_LOW_PREP_HIGH if the high cells have been sampled.
	localparam FSM_BITS = clogb2(5);
	localparam [FSM_BITS-1:0] RESET = 0;						  //% SST=0, WRSTRB=0, WR=X.
	localparam [FSM_BITS-1:0] RESET_WAIT = 1;               //% SST=0, WRSTRB=0, WR=X.
	localparam [FSM_BITS-1:0] SAMPLE_LOW_PREP_HIGH 		= 2; //% SST=1, WRSTRB=0, WR=HIGHBLOCK.
	localparam [FSM_BITS-1:0] SAMPLE_LOW_TRANSFER_HIGH = 3; //% SST=1, WRSTRB=1, WR=HIGHBLOCK.
	localparam [FSM_BITS-1:0] PREP_LOW_SAMPLE_HIGH		= 4; //% SST=0, WRSTRB=0, WR=LOWBLOCK.
	localparam [FSM_BITS-1:0] TRANSFER_LOW_SAMPLE_HIGH = 5; //% SST=0, WRSTRB=1, WR=LOWBLOCK.
	reg [FSM_BITS-1:0] state = RESET;							  //% State variable.
	assign dbg_state_o = state;
	
	//% Synchronization flop for SSp
	reg ssp_sync = 0;
	//% Copy of SSp sync for SSt
	reg sst_sync = 0;
	//% Synchronization flop for WRSTRB
	reg wrstrb_sync = 0;
	//% Acknowledge that a block has been written.
	reg wr_ack = 0;
	
	//% 1 if the high cells have been sampled to, 0 otherwise. (Used after reset).
	reg high_cells_sampled = 0;
	//% 1 if the low cells have been sampled to, 0 otherwise. Unused, here for completeness.
	reg low_cells_sampled = 0;
	//% Registered to ssp_sync on the next SSp rising edge, and sst_sync on the next clk_i edge.
	//% SSp/Sst go high on 2nd rising clock edge after ss_enable is true.
	wire ss_enable = (state == RESET && !rst_i) || (state == RESET_WAIT) || (state == PREP_LOW_SAMPLE_HIGH || state == TRANSFER_LOW_SAMPLE_HIGH);
	//% Registered to wrstrb_sync on next wrstrb clock rising edge. 
	//% WRSTRB goes high on 2nd rising clock edge after wrstrb_enable is true.
	wire wrstrb_enable = (state == SAMPLE_LOW_TRANSFER_HIGH || state == TRANSFER_LOW_SAMPLE_HIGH);

	always @(posedge clk_i) begin : FSM_LOGIC
		if (rst_i) state <= RESET;
		else begin
			case (state)
				RESET: state <= RESET_WAIT;
				RESET_WAIT: state <= SAMPLE_LOW_PREP_HIGH;
				SAMPLE_LOW_PREP_HIGH: state <= SAMPLE_LOW_TRANSFER_HIGH;
				SAMPLE_LOW_TRANSFER_HIGH: state <= PREP_LOW_SAMPLE_HIGH;
				PREP_LOW_SAMPLE_HIGH: state <= TRANSFER_LOW_SAMPLE_HIGH;
				TRANSFER_LOW_SAMPLE_HIGH: state <= SAMPLE_LOW_PREP_HIGH;
			endcase
		end
	end

	//% Acknowledge.
	always @(posedge clk_i) begin : ACK_LOGIC
		if (wr_ack) wr_ack <= 0;
		else if (((state == SAMPLE_LOW_PREP_HIGH && high_cells_sampled) || state == PREP_LOW_SAMPLE_HIGH) && enable_i) wr_ack <= 1;
	end

	//% High/low cell sampling indicator logic.
	always @(posedge clk_i) begin : CELLS_SAMPLED_LOGIC
		if (rst_i) begin
			high_cells_sampled <= 0;
			low_cells_sampled <= 0;
		end else begin
			if (state == SAMPLE_LOW_TRANSFER_HIGH) low_cells_sampled <= 1;
			if (state == TRANSFER_LOW_SAMPLE_HIGH) high_cells_sampled <= 1;
		end
	end

	//% Synchronization of SSp to ssp_clk domain
	always @(posedge clk_i) begin : SSP_SYNC_LOGIC
		ssp_sync <= ss_enable;
	end

	//% Copy of SSp sync for SSt.
	always @(posedge clk_i) begin : SST_SYNC_LOGIC
		sst_sync <= ss_enable;
	end

	//% Synchronization for WRSTRB.
	always @(posedge clk_i) begin : WRSTRB_SYNC_LOGIC
		wrstrb_sync <= wrstrb_enable;
	end

	//% Enable the latching of the write address. 1 cycle before PREP stages, so WR stable in PREP.
	wire latch_wr_address = (state == SAMPLE_LOW_TRANSFER_HIGH || state == TRANSFER_LOW_SAMPLE_HIGH);

	// Registers.
	generate
		genvar i;
		for (i=0;i<9;i=i+1) begin : WRFF
			// Write address registers.
			(* IOBUF = "TRUE" *) (* INIT = 0 *) FDE wr_ff(.D(wr_block_i[i]),.C(clk_i),.CE(latch_wr_address),.Q(wr_o[i]));
			// Debug write address registers.
			(* INIT = 0 *) FDE dbg_wr_ff(.D(wr_block_i[i]),.C(clk_i),.CE(latch_wr_address),.Q(dbg_wr_o[i]));
		end
		// WR[9] register
		(* IOBUF = "TRUE" *) (* INIT = 0 *) FDE wren_ff(.D(enable_i),.C(clk_i),.CE(latch_wr_address),.Q(wr_o[9]));
		// Debug WR[9] register
		(* INIT = 0 *) FDE dbg_wren_ff(.D(enable_i),.C(clk_i),.CE(latch_wr_address),.Q(dbg_wr_o[9]));
		// SSp register.
		(* IOBUF = "TRUE" *) (* INIT = 0 *) FDE ssp_ff(.D(ssp_sync),.C(ssp_clk_i),.CE(1'b1),.Q(ssp_o));
		// SSt register
		(* IOBUF = "TRUE" *) (* INIT = 0 *) FDE sst_ff(.D(sst_sync),.C(clk_i),.CE(1'b1),.Q(sst_o));
		// Debug versions of SSp, SSt register.
		(* INIT = 0 *) FDE dbg_ss_ff(.D(sst_sync),.C(clk_i),.CE(1'b1),.Q(dbg_sst_o));

		(* IOBUF = "TRUE" *) (* INIT = 0 *) FDE wrstrb_ff(.D(wrstrb_sync),.C(wrstrb_clk_i),.CE(1'b1),.Q(wrstrb_o));
		// Debug WRSTRB register
		(* INIT = 0 *) FDE dbg_wrstrb_ff(.D(wrstrb_sync),.C(clk_i),.CE(1'b1),.Q(dbg_wrstrb_o));
	endgenerate
	
	assign dbg_ssp_o = dbg_sst_o;
	assign wr_phase_o = ((state == SAMPLE_LOW_PREP_HIGH && high_cells_sampled) ||
								(state == TRANSFER_LOW_SAMPLE_HIGH));
	assign wr_ack_o = wr_ack;
endmodule

