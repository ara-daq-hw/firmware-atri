`timescale 1ns / 1ps
// IRS soft trigger control.
module irs_softtrig_ctrl(
		input [7:0] dat_i,
		output [7:0] dat_o,
		input wr_i,
		input clk_i,
		output trig_o
    );


endmodule
